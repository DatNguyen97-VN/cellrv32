// ##################################################################################################
// # << CELLRV32 - Processor-internal instruction memory (IMEM) >>                                  #
// # ********************************************************************************************** #
// # This memory optionally includes the in-place executable image of the application. See the      #
// # processor's documentary to get more information.                                               #
// # ********************************************************************************************** #
`ifndef  _INCL_DEFINITIONS
  `define _INCL_DEFINITIONS
  `include "cellrv32_package.svh"
`endif // _INCL_DEFINITIONS

// this package is generated by the image generator
import cellrv32_bootloader_image::*;

module cellrv32_boot_rom #(
    parameter logic [31:0] BOOTROM_BASE = 32'h00000000 // boot ROM base address
) (
    input  logic         clk_i,  // global clock line
    input  logic         rden_i, // read enable
    input  logic         wren_i, // write enable
    input  logic [31:0]  addr_i, // address
    output logic [31:0]  data_o, // data out
    output logic         ack_o,  // transfer acknowledge
    output logic         err_o   // transfer error
);
    /* determine required ROM size in bytes (expand to next power of two) */
    localparam int boot_rom_size_index_c = index_size_f($size(bootloader_init_image)); // address with (32-bit entries)
    localparam int boot_rom_size_c       = (2**boot_rom_size_index_c)*4; // size in bytes

    /* IO space: module base address */
    localparam int hi_abb_c = 31; // high address boundary bit
    localparam int lo_abb_c = index_size_f(boot_rom_max_size_c); // low address boundary bit
    
    /* local signals */
    logic acc_en;
    logic rden;
    logic [31:0] rdata;
    logic [boot_rom_size_index_c-1:0] addr;

    /* ROM - initialized with executable code */
    const logic [31:0] mem_rom [16*1024] = mem32_init_boot_f(bootloader_init_image, boot_rom_max_size_c/4);

    // Sanity Checks -----------------------------------------------------------------------------
    // -------------------------------------------------------------------------------------------
    initial begin
        assert (1'b0) else $info("CELLRV32 PROCESSOR CONFIG NOTE: Implementing internal bootloader ROM (%0d bytes)", boot_rom_size_c);
        assert (boot_rom_size_c <= boot_rom_max_size_c) else $error("CELLRV32 PROCESSOR CONFIG ERROR! Boot ROM size out of range! Max %0d bytes", boot_rom_max_size_c);
    end

    // Access Control ----------------------------------------------------------------------------
    // -------------------------------------------------------------------------------------------
    assign acc_en = (addr_i[hi_abb_c : lo_abb_c] == BOOTROM_BASE[hi_abb_c : lo_abb_c]) ? 1'b1 : 1'b0;
    assign addr   = addr_i[boot_rom_size_index_c+1 : 2]; // word aligned

    // Memory Access -----------------------------------------------------------------------------
    // -------------------------------------------------------------------------------------------
    always_ff @( posedge clk_i ) begin : mem_file_access
      rden  <= acc_en & rden_i;
      err_o <= acc_en & wren_i;
      // reduce switching activity when not accessed
      if (acc_en) begin
        rdata <= mem_rom[addr];
      end
    end : mem_file_access

    /* output gate */
    assign data_o = rden ? rdata : '0;
    assign ack_o = rden;

endmodule